module input_reg
  (
  in
  );

input [15:0] in;

parameter REG = 0;// Marks this module as a register
parameter ADDR = 0; // Address of register

endmodule
